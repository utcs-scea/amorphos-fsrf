// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

// Used with modifications by Joshua Landgraf

`ifndef CL_DRAM_DMA_PKG
`define CL_DRAM_DMA_PKG
 
interface axi_bus_t;
   logic[15:0] awid;
   logic[63:0] awaddr;
   logic[7:0] awlen;
   logic[2:0] awsize;
   logic awvalid;
   logic awready;
   
   logic[511:0] wdata;
   logic[63:0] wstrb;
   logic wlast;
   logic wuser;
   logic wvalid;
   logic wready;
   
   logic[15:0] bid;
   logic[1:0] bresp;
   logic bvalid;
   logic bready;
   
   logic[15:0] arid;
   logic[63:0] araddr;
   logic[7:0] arlen;
   logic[2:0] arsize;
   logic arvalid;
   logic arready;
   
   logic[15:0] rid;
   logic[511:0] rdata;
   logic[1:0] rresp;
   logic ruser;
   logic rlast;
   logic rvalid;
   logic rready;

   modport master (input awid, awaddr, awlen, awsize, awvalid, output awready,
                  input wdata, wstrb, wlast, wuser, wvalid, output wready,
                  output bid, bresp, bvalid, input bready,
                  input arid, araddr, arlen, arsize, arvalid, output arready,
                  output rid, rdata, rresp, rlast, ruser, rvalid, input rready);

   modport slave (output awid, awaddr, awlen, awsize, awvalid, input awready,
                  output wdata, wstrb, wlast, wuser, wvalid, input wready,
                  input bid, bresp, bvalid, output bready,
                  output arid, araddr, arlen, arsize, arvalid, input arready,
                  input rid, rdata, rresp, rlast, ruser, rvalid, output rready);
endinterface

`endif //CL_DRAM_DMA_PKG
