`define max_layers 3
`define num_pe 4
`define num_pu 1

`define max_rd_mem_idx 3
`define max_wr_mem_idx 3
