`ifndef USER_PARAMS_SV_INCLUDED
`define USER_PARAMS_SV_INCLUDED
                        
package UserParams;

parameter NUM_APPS = 4;
parameter CONFIG_APPS = 10;

endpackage
`endif 
